package env_pack;
   import uvm_pkg::*;
   import agent_pack::*;
`include "uvm_macros.svh"
`include "Scoreboard.svh"
`include "env_config.svh"
`include "Environment.svh"
endpackage // env_pack
   