package agent_pack;
   import uvm_pkg::*
`include "uvm_macros.svh"
`include "Transaction.svh"
`include "Sequence.svh"
`include "Sequencer.svh"
`include "Driver.svh"
`include "Monitor.svh"
`include "agent_config.svh"
`include "Agent.svh"

endpackage // agent_pack
   