package test_pack ;
   import uvm_pkg::*;
   import env_pack::*;
`include "uvm_macros.svh"
`include "test.svh"
endpackage // test_pack
   